

https://edaplayground.com/x/Wxqr

https://edaplayground.com/x/gvh_
